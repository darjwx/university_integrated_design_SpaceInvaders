----------------------------------------------------------------------------------
-- Company: UC3M
-- Engineers: Dario Jimenez Juiz
--            Gabriel Minelli Lli
--            Alvaro Manzanero Moran
--
-- Create Date: 07.10.2019 11:44:18
-- Module Name: formatoVGA - Behavioral
-- Project Name: SpaceInv
-- Description: Definicion y control de lo que se muestra por pantalla.
--              Ligado al bloque vga.
--
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.NUMERIC_STD.all;

entity formatoVGA is
    Port ( X : in UNSIGNED (9 downto 0);
           Y : in UNSIGNED (9 downto 0);
           test : in std_logic;
           invadersH : in unsigned (0 to 19);
           invadersV : in integer range 0 to 14;
           naveH : in integer range 0 to 19;
           disparoH : in integer range 0 to 19;
           disparoV : in integer range 0 to 14;
           mensajeV : in std_logic;
           mensajeD : in std_logic;
           Color : out UNSIGNED (2 downto 0));
end formatoVGA;

architecture Behavioral of formatoVGA is
--Señales que contienen la parte alta o baja de las señales de entrada X,Y
signal rX: integer range 0 to 19;
signal rY: integer range 0 to 14;
signal detailX: integer range 0 to 31;
signal detailY: integer range 0 to 31;

--Señales que contienen la parte alta o baja de X,Y en formato de entero
signal upX : unsigned (4 downto 0);
signal upY : unsigned (4 downto 0);
signal downX: unsigned (4 downto 0);
signal downY: unsigned (4 downto 0);


-- Matriz 32*32
type icono is array (0 to 31, 0 to 31) of std_logic;

--Icono que se mostrara cuando el jugador gane
constant victoria : icono := ("00100000000000000000000000000100",
                              "00010000000000000000000000001000",
                              "00001000000000000000000000010000",
                              "00000100000000000000000000100000",
                              "00000010000000000000000001000000",
                              "00000001000000000000000010000000",
                              "00000000100000000000000100000000",
                              "00000000010000000000001000000000",
                              "00000000001000000000010000000000",
                              "00000000000100000000100000000000",
                              "00000000000010000001000000000000",
                              "00000000000001000010000000000000",
                              "00000000000000100100000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000000000000000000000",
                              "00000000000000000000000000000000",
                              "00000000000000000000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000",
                              "00000000000000011000000000000000");

--Icono que se mostrara cuando el jugador sea derrotado
constant derrota : icono := ( "11110000000000000000000000000000",
                              "11001100000000000000000000000000",
                              "11000011000000000000000000000000",
                              "11000000110000000000000000000000",
                              "11000000001100000000000000000000",
                              "11000000000011000000000000000000",
                              "11000000000000110000000000000000",
                              "11000000000000001100000000000000",
                              "11000000000000000011000000000000",
                              "11000000000000000000110000000000",
                              "11000000000000000000001100000000",
                              "11000000000000000000000011000000",
                              "11000000000000000000000000110000",
                              "11000000000000000000000000001100",
                              "11000000000000000000000000001100",
                              "11000000000000000000000000110000",
                              "11000000000000000000000011000000",
                              "11000000000000000000001100000000",
                              "11000000000000000000110000000000",
                              "11000000000000000011000000000000",
                              "11000000000000011000000000000000",
                              "11000000000001100000000000000000",
                              "11000000000110000000000000000000",
                              "11000000011000000000000000000000",
                              "11000001100000000000000000000000",
                              "11000110000000000000000000000000",
                              "11111000000000000000000000000000",
                              "11111111111100000000000000000000",
                              "11000000000000000000000000000000",
                              "11111111111100000000000000000000",
                              "11000000000000000000000000000000",
                              "11111111111100000000000000000000");

--Icono que representa a los invasorres
constant invasores : icono := ("00111100000000000000000000111100",
                               "00111100000000000000000000111100",
                               "00111100000000000000000000111100",
                               "00111100000000000000000000111100",
                               "00000011110000000000001111000000",
                               "00000011110000000000001111000000",
                               "00000011110000000000001111000000",
                               "00000011110000000000001111000000",
                               "00111111111111111111111111111100",
                               "00111111111111111111111111111100",
                               "00111111111111111111111111111100",
                               "00111111111111111111111111111100",
                               "00111100001111111111110000111100",
                               "00111100001111111111110000111100",
                               "00111100001111111111110000111100",
                               "00111100001111111111110000111100",
                               "00111111111111111111111111111100",
                               "00111111111111111111111111111100",
                               "00111111111111111111111111111100",
                               "00111111111111111111111111111100",
                               "00111111111111111111111111111100",
                               "00111111111111111111111111111100",
                               "00111111111111111111111111111100",
                               "00111111111111111111111111111100",
                               "00111100000000000000000000111100",
                               "00111100000000000000000000111100",
                               "00111100000000000000000000111100",
                               "00111100000000000000000000111100",
                               "00000011111111000011111111000000",
                               "00000011111111000011111111000000",
                               "00000011111111000011111111000000",
                               "00000011111111000011111111000000");

--Icono que representa a la bala
constant bala : icono := ("00000000000000000000000000000000",
                          "00000000000000000000000000000000",
                          "00000000000000000000000000000000",
                          "00000000000000000000000000000000",
                          "00000000000000000000000000000000",
                          "00000000000000000000000000000000",
                          "00000000000000000000000000000000",
                          "00000000000000000000000000000000",
                          "00000000000000011000000000000000",
                          "00000000000000011000000000000000",
                          "00000000000000011000000000000000",
                          "00000000000000011000000000000000",
                          "00000000000000011000000000000000",
                          "00000000000000011000000000000000",
                          "00000000000000011000000000000000",
                          "00000000000000011000000000000000",
                          "00000000000000111100000000000000",
                          "00000000000000111000000000000000",
                          "00000000000000111100000000000000",
                          "00000000000000111100000000000000",
                          "00000000000000111100000000000000",
                          "00000000000001111110000000000000",
                          "00000000000011111111000000000000",
                          "00000000001111111111110000000000",
                          "00000000000010011001000000000000",
                          "00000000000001010010000000000000",
                          "00000000000000101000000000000000",
                          "00000000000000010000000000000000",
                          "00000000000000000000000000000000",
                          "00000000000000000000000000000000",
                          "00000000000000000000000000000000",
                          "00000000000000000000000000000000");

--Icono que representa a la nave
constant nave : icono := ("00000000000000111100000000000000",
                          "00000000000000111100000000000000",
                          "00000000000000111100000000000000",
                          "00000000000000111100000000000000",
                          "00000000000000111100000000000000",
                          "00000000000000111100000000000000",
                          "00110000001111111111110000001100",
                          "00110000001111111111110000001100",
                          "00110000001111111111110000001100",
                          "00110000001111111111110000001100",
                          "00110000111111111111111100001100",
                          "00110000111111111111111100001100",
                          "11111111111111111111111111111111",
                          "11111111111111111111111111111111",
                          "11111111111111111111111111111111",
                          "11111111111111111111111111111111",
                          "11111111111111111111111111111111",
                          "11111111111111111111111111111111",
                          "11111111111111111111111111111111",
                          "11111111111111111111111111111111",
                          "11111111111111111111111111111111",
                          "11111111111111111111111111111111",
                          "11110000111111111111111100001111",
                          "11110000111111111111111100001111",
                          "11110000001111111111110000001111",
                          "11110000001111111111110000001111",
                          "00000000001100000000110000000000",
                          "00000000001100000000110000000000",
                          "00000000110000000000001100000000",
                          "00000000110000000000001100000000",
                          "00000000110000000000001100000000",
                          "00000000110000000000001100000000");





begin


-- Warning Y(9) not connected
-- 5 bits > que lo que puede almacenar rY (integer 0 to 14)
  upX <= X(9)&X(8)&X(7)&X(6)&X(5);
  upY <= Y(9)&Y(8)&Y(7)&Y(6)&Y(5);
  downX <= X(4)&X(3)&X(2)&X(1)&X(0);
  downY <= Y(4)&Y(3)&Y(2)&Y(1)&Y(0);

  --Transforma la parte alta o baja de X,Y en enteros
  process(upX,upY,downX,downY)
  begin
    rX <= to_integer(upX);
    rY <= to_integer(upY);
    detailX <= to_integer(downX);
    detailY <= to_integer(downY);
  end process;

 --Define la imagen que se va a mostrar por pantalla y sus colores
 process(rX,rY,test,invadersH,invadersV,upX,upY,naveH,disparoH,disparoV,mensajeV,mensajeD,detailX,detailY)
 begin
   if test = '0' then
     --Mensaje de victoria
     if mensajeV = '1' then
        if victoria(detailY,detailX) = '1' then
          Color <= "010";
        else
          Color <= "000";
        end if;
     --Mensaje de derrota
     elsif mensajeD = '1' then
       if derrota(detailY,detailX) = '1' then
         Color <= "100";
       else
         Color <= "000";
       end if;
     elsif rX <= 19 and rY <= 14 then
         --Invasores
         if invadersH(rX) = '1' and rY = invadersV then
           if invasores(detailY,detailX) = '1' then
             Color <= "010";
           else
             Color <= "000";
           end if;
         elsif rX = naveH and rY = 14 then
           --Nave
           if nave(detailY,detailX) = '1' then
             Color <= "110";
           else
             Color <= "000";
           end if;
         elsif rX = disparoH and rY = disparoV then
           --Bala
           if bala(detailY,detailX) = '1' then
             Color <= "100";
           else
             Color <= "000";
           end if;
         else
           Color <= "000";
         end if;
     else
       Color <= "000";
     end if;
   else
     --Tablero
       if (upX(0) = '1' and upY(0) = '1') or (upX(0) = '0' and upY(0) = '0') then
         -- Blanco
         Color <= "111";
       else
         -- Negro
         Color <= "000";
       end if;
     end if;
 end process;


end Behavioral;
